module alu (
    input wire                 clk_in;
    input wire                 rst_in;
    input wire                 rdy_in;

    input wire                 opType;

    output reg                 aluResult;
);

always @(posedge clk_in) begin

end