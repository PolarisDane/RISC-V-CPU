module rob (
    input wire                      clk_in,
    input wire                      rst_in,
    input wire                      rdy_in,

    input wire                      dc_to_rob,
    output reg                      rob_to_if_alter_pc,
    output reg                      rob_to_if_alter_pc_ready,
)
endmodule