module InstructionUnit (
    
);