module lsb (
    input wire                      clk_in,
    input wire                      rst_in,
    input wire                      rdy_in,

    input wire                      dc_to_lsb_,




    input wire                      mc_to_lsb_
    output reg                      lsb_to_mc_ready,
    output reg                      lsb_to_mc_op,
    output reg                      lsb_to_mc_opType,
    output reg                      lsb_to_mc_
)

endmodule